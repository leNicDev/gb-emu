module ppu

pub fn init() {

}

pub fn tick() {
	
}