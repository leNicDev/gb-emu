module timer

pub fn init() {

}

pub fn tick() {
	
}